`timescale 1ns/1ps

module mux_tb;

reg [31:0] I0;
reg [31:0] I1;
reg [31:0] I2;
reg [31:0] I3;
reg [1:0] S;

wire [31:0] Y;

MUX32_4x1 mux_4x1inst(.Y(Y), .I0(I0), .I1(I1), .I2(I2), .I3(I3), .S(S));
initial
begin
#5 I0='b1111; I1='b1010; I2='b0001; I3='b0000; S='b00;

#5 I0='b1111; I1='b1010; I2='b0001; I3='b0000; S='b10;
#5 I0='b1111; I1='b1010; I2='b0001; I3='b0000; S='b01;
#5 I0='b1111; I1='b1010; I2='b0001; I3='b0000; S='b11;
#5;
end


reg [31:0] I4;
reg [31:0] I5;
reg [31:0] I6;
reg [31:0] I7;
reg [2:0] Q;
wire [31:0] R;

MUX32_8x1 mux_8x1inst(.Y(R), .I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .I6(I6), .I7(I7),.S(Q));
initial
begin
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b000;
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b001;
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b010;
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b011;
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b100;
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b101;
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b110;
#5 I0='b0000; I1='b0001; I2='b0010; I3='b0011; I4='b0100; I5='b0101; I6='b0110; I7='b0111; Q='b111;
#5;
end

reg [31:0] R0;
reg [31:0] R1;
reg [31:0] R2;
reg [31:0] R3;
reg [31:0] R4;
reg [31:0] R5;
reg [31:0] R6;
reg [31:0] R7;
reg [31:0] R8;
reg [31:0] R9;
reg [31:0] R10;
reg [31:0] R11;
reg [31:0] R12;
reg [31:0] R13;
reg [31:0] R14;
reg [31:0] R15;
reg [3:0] M;
wire [31:0] B;

MUX32_16x1 mux_16x1(.Y(B), .I0(R0), .I1(R1), .I2(R2), .I3(R3), .I4(R4), .I5(R5), .I6(R6), .I7(R7),
                     .I8(R8), .I9(R9), .I10(R10), .I11(R11), .I12(R12), .I13(R13), .I14(R14), .I15(R15), .S(M));
initial
begin
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0000;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0001;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0010;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0011;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0100;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0101;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0110;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b0111;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1000;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1001;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1010;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1011;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1100;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1101;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1110;
#5 R0='b00000; R1='b00001; R2='b00010; R3='b00011; R4='b00100; R5='b00101; R6='b00110; R7='b00111;
	R8='b01000; R9='b01001; R10='b01010; R11='b01011; R12='b01100; R13='b01101; R14='b01111; R15='b10000; M='b1111;
#5;
end

endmodule